library verilog;
use verilog.vl_types.all;
entity Register8_vlg_vec_tst is
end Register8_vlg_vec_tst;
