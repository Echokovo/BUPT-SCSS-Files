library verilog;
use verilog.vl_types.all;
entity Encoder8421toGray_vlg_vec_tst is
end Encoder8421toGray_vlg_vec_tst;
