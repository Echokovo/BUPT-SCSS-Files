library verilog;
use verilog.vl_types.all;
entity Decoder3to8_vlg_vec_tst is
end Decoder3to8_vlg_vec_tst;
