library verilog;
use verilog.vl_types.all;
entity compare4_vlg_vec_tst is
end compare4_vlg_vec_tst;
