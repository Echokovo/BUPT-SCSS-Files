library verilog;
use verilog.vl_types.all;
entity String_Detector_vlg_vec_tst is
end String_Detector_vlg_vec_tst;
