library verilog;
use verilog.vl_types.all;
entity compare4_vlg_check_tst is
    port(
        YA              : in     vl_logic;
        YB              : in     vl_logic;
        YC              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end compare4_vlg_check_tst;
