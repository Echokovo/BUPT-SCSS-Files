library verilog;
use verilog.vl_types.all;
entity Count4_vlg_vec_tst is
end Count4_vlg_vec_tst;
