library verilog;
use verilog.vl_types.all;
entity Fulladder_vlg_vec_tst is
end Fulladder_vlg_vec_tst;
